module vglyph

import gg
import math

// hit_test_rect returns the bounding box of the character at (x, y) relative to the layout origin.
// Returns none if no character is found close enough.
pub fn (l Layout) hit_test_rect(x f32, y f32) ?gg.Rect {
	for cr in l.char_rects {
		if x >= cr.rect.x && x <= cr.rect.x + cr.rect.width && y >= cr.rect.y
			&& y <= cr.rect.y + cr.rect.height {
			return cr.rect
		}
	}
	return none
}

// get_char_rect returns the bounding box for a specific character byte index.
pub fn (l Layout) get_char_rect(index int) ?gg.Rect {
	rect_idx := l.char_rect_by_index[index] or { return none }
	return l.char_rects[rect_idx].rect
}

// hit_test returns the byte index of the character at (x, y) relative to origin.
// Returns -1 if no character is found.
//
// Algorithm:
// Linear search (O(N)) over baked char rects.
// Trade-offs:
// - Efficiency: Faster than spatial structures for typical N < 1000.
// - Accuracy: Returns first matching index (logical order).
pub fn (l Layout) hit_test(x f32, y f32) int {
	// Simple linear search.
	// We could optimize with spatial partitioning if needed.
	for cr in l.char_rects {
		if x >= cr.rect.x && x <= cr.rect.x + cr.rect.width && y >= cr.rect.y
			&& y <= cr.rect.y + cr.rect.height {
			return cr.index
		}
	}
	return -1
}

// get_closest_offset returns the byte index of the character closest to (x, y).
// Handles clicks outside bounds (returns nearest edge/line).
pub fn (l Layout) get_closest_offset(x f32, y f32) int {
	if l.lines.len == 0 {
		return 0
	}

	// 1. Find the closest line vertically
	mut closest_line_idx := 0
	mut min_dist_y := f32(1e9)

	for i, line in l.lines {
		// Check containment or distance
		// Simple distance to vertical center of line
		line_mid_y := line.rect.y + line.rect.height / 2
		dist := match true {
			y >= line.rect.y && y <= line.rect.y + line.rect.height { 0.0 } // Inside
			else { math.abs(y - line_mid_y) }
		}

		if dist < min_dist_y {
			min_dist_y = dist
			closest_line_idx = i
		}
	}

	target_line := l.lines[closest_line_idx]

	// 2. Resolve X using Pango (requires recalculation or stored PangoLayout... wait)
	// We don't have the PangoLayout stored in V struct Layout (it's transient).
	// So we must rely on our cached data (CharRects).

	// Linear search within the line's range
	line_end := target_line.start_index + target_line.length
	mut closest_char_idx := target_line.start_index
	mut min_dist_x := f32(1e9)

	// If x is before line start
	if x < target_line.rect.x {
		return target_line.start_index
	}
	// If x is after line end
	if x > target_line.rect.x + target_line.rect.width {
		// Return end of line (but we need to know if it's newline char or not)
		// Usually target_line.start_index + target_line.length
		return line_end
	}

	// Scan chars in this line using O(1) index lookup
	for i in target_line.start_index .. line_end {
		rect_idx := l.char_rect_by_index[i] or { continue }
		cr := l.char_rects[rect_idx]
		char_mid_x := cr.rect.x + cr.rect.width / 2
		dist := math.abs(x - char_mid_x)
		if dist < min_dist_x {
			min_dist_x = dist
			closest_char_idx = i
		}
	}

	// Edge case: if we are closer to the right edge of the last char
	// we should probably return index + char_len?
	// Simplified: return index of char center closest to mouse.
	return closest_char_idx
}

// get_selection_rects returns a list of rectangles covering the text range [start, end).
pub fn (l Layout) get_selection_rects(start int, end int) []gg.Rect {
	if start >= end || l.lines.len == 0 {
		return []gg.Rect{}
	}

	mut rects := []gg.Rect{}
	mut s := start
	mut e := end

	// Clamp
	if s < 0 {
		s = 0
	}
	// Max index? approximation
	// if e > max_len { ... }

	for line in l.lines {
		line_end := line.start_index + line.length

		// Check intersection
		// Range 1: [line.start, line_end)
		// Range 2: [s, e)

		overlap_start := if s > line.start_index { s } else { line.start_index }
		overlap_end := if e < line_end { e } else { line_end }

		if overlap_start < overlap_end {
			// Calculate visual rect for this overlap using O(1) index lookup
			mut min_x := f32(1e9)
			mut max_x := f32(-1e9)
			mut found := false

			for i in overlap_start .. overlap_end {
				rect_idx := l.char_rect_by_index[i] or { continue }
				cr := l.char_rects[rect_idx]
				if cr.rect.x < min_x {
					min_x = cr.rect.x
				}
				if cr.rect.x + cr.rect.width > max_x {
					max_x = cr.rect.x + cr.rect.width
				}
				found = true
			}

			if found {
				rects << gg.Rect{
					x:      min_x
					y:      line.rect.y
					width:  max_x - min_x
					height: line.rect.height
				}
			}
		}
	}
	return rects
}

// get_font_name_at_index returns the family name of the font used to render
// the character at the given byte index.
pub fn (l Layout) get_font_name_at_index(index int) string {
	for item in l.items {
		if index >= item.start_index && index < item.start_index + item.length {
			if item.ft_face != unsafe { nil } {
				return unsafe { cstring_to_vstring(item.ft_face.family_name) }
			}
		}
	}
	return 'Unknown'
}

// get_cursor_pos returns the geometry for rendering a cursor at the given byte index.
// Returns none if index is out of bounds.
//
// Algorithm:
// 1. Check bounds (0 <= byte_index <= text length via log_attrs.len - 1)
// 2. Try exact char_rect lookup for index
// 3. If at line end, use line rect right edge
// 4. Return x (left edge of char or line end), y (line top), height (line height)
//
// Note: This uses cached char_rects/lines. For precise bidi cursor positioning,
// a future version could store cursor_pos during layout build from Pango.
pub fn (l Layout) get_cursor_pos(byte_index int) ?CursorPosition {
	// Bounds check using log_attrs (len = text_len + 1)
	if l.log_attrs.len == 0 {
		return none
	}
	max_index := l.log_attrs.len - 1
	if byte_index < 0 || byte_index > max_index {
		return none
	}

	// Try exact char rect lookup
	if rect := l.get_char_rect(byte_index) {
		return CursorPosition{
			x:      rect.x
			y:      rect.y
			height: rect.height
		}
	}

	// Fallback: find containing line
	for line in l.lines {
		line_end := line.start_index + line.length
		if byte_index >= line.start_index && byte_index <= line_end {
			if byte_index == line_end {
				// At end of line - cursor at right edge
				return CursorPosition{
					x:      line.rect.x + line.rect.width
					y:      line.rect.y
					height: line.rect.height
				}
			}
			// At start of line
			return CursorPosition{
				x:      line.rect.x
				y:      line.rect.y
				height: line.rect.height
			}
		}
	}

	// Ultimate fallback: use first line if exists
	if l.lines.len > 0 {
		first_line := l.lines[0]
		return CursorPosition{
			x:      first_line.rect.x
			y:      first_line.rect.y
			height: first_line.rect.height
		}
	}

	return none
}

// move_cursor_left returns the byte index of the previous valid cursor position.
// Returns current index if already at start. Respects grapheme clusters (won't land inside emoji).
pub fn (l Layout) move_cursor_left(byte_index int) int {
	if byte_index <= 0 || l.log_attrs.len == 0 {
		return 0
	}
	// Scan backwards for previous is_cursor_position
	for i := byte_index - 1; i >= 0; i-- {
		if i < l.log_attrs.len && l.log_attrs[i].is_cursor_position {
			return i
		}
	}
	return 0
}

// move_cursor_right returns the byte index of the next valid cursor position.
// Returns current index if already at end. Respects grapheme clusters.
pub fn (l Layout) move_cursor_right(byte_index int) int {
	if l.log_attrs.len == 0 {
		return byte_index
	}
	max_index := l.log_attrs.len - 1
	if byte_index >= max_index {
		return max_index
	}
	// Scan forward for next is_cursor_position
	for i in (byte_index + 1) .. l.log_attrs.len {
		if l.log_attrs[i].is_cursor_position {
			return i
		}
	}
	return max_index
}

// move_cursor_word_left returns the byte index of the previous word start.
// Skips to word boundary, not just cursor position.
pub fn (l Layout) move_cursor_word_left(byte_index int) int {
	if byte_index <= 0 || l.log_attrs.len == 0 {
		return 0
	}
	// First move left to skip current position
	mut idx := byte_index - 1
	// Skip any whitespace/non-word chars
	for idx > 0 && !l.log_attrs[idx].is_word_start {
		idx--
	}
	// If we found a word start, return it
	if idx >= 0 && l.log_attrs[idx].is_word_start {
		return idx
	}
	return 0
}

// move_cursor_word_right returns the byte index of the next word start.
pub fn (l Layout) move_cursor_word_right(byte_index int) int {
	if l.log_attrs.len == 0 {
		return byte_index
	}
	max_index := l.log_attrs.len - 1
	if byte_index >= max_index {
		return max_index
	}
	// Scan forward for next word start
	for i in (byte_index + 1) .. l.log_attrs.len {
		if l.log_attrs[i].is_word_start {
			return i
		}
	}
	return max_index
}

// move_cursor_line_start returns the byte index of the start of the current line.
pub fn (l Layout) move_cursor_line_start(byte_index int) int {
	for line in l.lines {
		line_end := line.start_index + line.length
		if byte_index >= line.start_index && byte_index <= line_end {
			return line.start_index
		}
	}
	// Fallback: return 0
	return 0
}

// move_cursor_line_end returns the byte index of the end of the current line.
pub fn (l Layout) move_cursor_line_end(byte_index int) int {
	for line in l.lines {
		line_end := line.start_index + line.length
		if byte_index >= line.start_index && byte_index <= line_end {
			return line_end
		}
	}
	// Fallback: return max index
	if l.log_attrs.len > 0 {
		return l.log_attrs.len - 1
	}
	return 0
}

// move_cursor_up returns byte index on previous line at similar x position.
// preferred_x is the x coordinate to try to maintain (pass -1 to use cursor's current x).
pub fn (l Layout) move_cursor_up(byte_index int, preferred_x f32) int {
	if l.lines.len == 0 {
		return byte_index
	}

	// Find current line index
	mut current_line_idx := -1
	mut target_x := preferred_x
	for i, line in l.lines {
		line_end := line.start_index + line.length
		if byte_index >= line.start_index && byte_index <= line_end {
			current_line_idx = i
			// If no preferred_x, use current cursor x
			if target_x < 0 {
				if pos := l.get_cursor_pos(byte_index) {
					target_x = pos.x
				} else {
					target_x = line.rect.x
				}
			}
			break
		}
	}

	if current_line_idx <= 0 {
		// Already on first line or not found
		return byte_index
	}

	// Find closest char on previous line
	prev_line := l.lines[current_line_idx - 1]
	return l.find_closest_index_in_line(prev_line, target_x)
}

// move_cursor_down returns byte index on next line at similar x position.
pub fn (l Layout) move_cursor_down(byte_index int, preferred_x f32) int {
	if l.lines.len == 0 {
		return byte_index
	}

	// Find current line index
	mut current_line_idx := -1
	mut target_x := preferred_x
	for i, line in l.lines {
		line_end := line.start_index + line.length
		if byte_index >= line.start_index && byte_index <= line_end {
			current_line_idx = i
			if target_x < 0 {
				if pos := l.get_cursor_pos(byte_index) {
					target_x = pos.x
				} else {
					target_x = line.rect.x
				}
			}
			break
		}
	}

	if current_line_idx < 0 || current_line_idx >= l.lines.len - 1 {
		// Not found or already on last line
		return byte_index
	}

	// Find closest char on next line
	next_line := l.lines[current_line_idx + 1]
	return l.find_closest_index_in_line(next_line, target_x)
}

// find_closest_index_in_line returns the byte index closest to target_x within the given line.
fn (l Layout) find_closest_index_in_line(line Line, target_x f32) int {
	line_end := line.start_index + line.length
	mut closest_idx := line.start_index
	mut min_dist := f32(1e9)

	for i in line.start_index .. line_end {
		rect_idx := l.char_rect_by_index[i] or { continue }
		cr := l.char_rects[rect_idx]
		char_mid_x := cr.rect.x + cr.rect.width / 2
		dist := math.abs(target_x - char_mid_x)
		if dist < min_dist {
			min_dist = dist
			closest_idx = i
		}
	}

	// Check if closer to end of line
	end_x := line.rect.x + line.rect.width
	if math.abs(target_x - end_x) < min_dist {
		return line_end
	}

	return closest_idx
}
