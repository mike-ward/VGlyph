module text_render

import gg
import time
import hash.fnv1a

struct CachedLayout {
mut:
	layout      Layout
	last_access i64
}

pub struct TextSystem {
mut:
	ctx          &Context
	renderer     &Renderer
	cache        map[u64]&CachedLayout
	eviction_age i64 = 5000 // ms
}

// new_text_system creates a new TextSystem.
// It initializes the underlying Pango context and the Renderer.
pub fn new_text_system(mut gg_ctx gg.Context) !&TextSystem {
	tr_ctx := new_context()!
	renderer := new_renderer(mut gg_ctx)
	return &TextSystem{
		ctx:      tr_ctx
		renderer: renderer
		cache:    map[u64]&CachedLayout{}
	}
}

// draw_text renders the given text string at coordinates (x, y) using the provided configuration.
// It automatically handles layout caching to optimize performance for repeated calls. [TextConfig](#TextConfig)
pub fn (mut ts TextSystem) draw_text(x f32, y f32, text string, cfg TextConfig) ! {
	key := ts.get_cache_key(text, cfg)
	ts.prune_cache()

	if key in ts.cache {
		mut item := ts.cache[key] or {
			return error('cache coherency error: key found but access failed')
		}
		item.last_access = time.ticks()
		ts.renderer.draw_layout(item.layout, x, y)
	} else {
		// Cache miss
		layout := ts.ctx.layout_text(text, cfg) or { return err }
		ts.cache[key] = &CachedLayout{
			layout:      layout
			last_access: time.ticks()
		}
		ts.renderer.draw_layout(layout, x, y)
	}
}

// text_width calculates and returns the width (in pixels) of the text if it were rendered with the given config.
// This is useful for layout calculations before rendering. [TextConfig](#TextConfig)
pub fn (mut ts TextSystem) text_width(text string, cfg TextConfig) !f32 {
	// For width we need the layout.
	// Difficult to guess without Pango shaping it.
	key := ts.get_cache_key(text, cfg)

	if key in ts.cache {
		mut item := ts.cache[key] or {
			return error('cache coherency error: key found but access failed')
		}
		item.last_access = time.ticks()
		return ts.get_layout_width(item.layout)
	}

	layout := ts.ctx.layout_text(text, cfg) or { return err }
	ts.cache[key] = &CachedLayout{
		layout:      layout
		last_access: time.ticks()
	}
	return ts.get_layout_width(layout)
}

// text_height calculates and returns the visual height (in pixels) of the text.
// This corresponds to the vertical space the text would occupy. [TextConfig](#TextConfig)
pub fn (mut ts TextSystem) text_height(text string, cfg TextConfig) !f32 {
	key := ts.get_cache_key(text, cfg)

	if key in ts.cache {
		mut item := ts.cache[key] or {
			return error('cache coherency error: key found but access failed')
		}
		item.last_access = time.ticks()
		return ts.renderer.max_visual_height(item.layout)
	}

	layout := ts.ctx.layout_text(text, cfg) or { return err }
	ts.cache[key] = &CachedLayout{
		layout:      layout
		last_access: time.ticks()
	}
	return ts.renderer.max_visual_height(layout)
}

// commit should be called at the end of the frame to upload the texture atlas.
pub fn (mut ts TextSystem) commit() {
	ts.renderer.commit()
}

// get_atlas_image returns the underlying texture atlas image.
// This is primarily for debugging purposes to visualize the safe-packing of glyphs.
pub fn (ts &TextSystem) get_atlas_image() gg.Image {
	return ts.renderer.atlas.image
}

// Internal Helpers

fn (ts TextSystem) get_cache_key(text string, cfg TextConfig) u64 {
	// Construct a unique key for the text + config combination
	// Format: text|font|width|align|wrap|markup|color|bg|u|s
	// Hash this string to get a compact u64 key
	s := '${text}|${cfg.font_name}|${cfg.width}|${cfg.align}|${cfg.wrap}|${cfg.use_markup}|${cfg.color}|${cfg.bg_color}|${cfg.underline}|${cfg.strikethrough}'
	return fnv1a.sum64_string(s)
}

fn (mut ts TextSystem) prune_cache() {
	now := time.ticks()

	if ts.cache.len < 100 {
		return
	}

	// simpler: usage of `keys()` copies the keys, so safe to delete.
	keys := ts.cache.keys()
	for k in keys {
		item := ts.cache[k] or { continue }
		if now - item.last_access > ts.eviction_age {
			ts.cache.delete(k)
		}
	}
}

fn (ts TextSystem) get_layout_width(layout Layout) f32 {
	// Layout width is usually the width of the widest line.
	// Pango layout already forced a width if wrapping, but if not wrapping, it'ss the max/sum of run widths.
	// `layout.items` has runs.
	mut max_x := f64(0)
	for item in layout.items {
		right := item.x + item.width
		if right > max_x {
			max_x = right
		}
	}
	return f32(max_x)
}
